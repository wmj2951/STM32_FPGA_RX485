module  lcd_char(
    input              sys_clk ,
    input              sys_rst_n ,
    //字符接口 
    input    [15:0]    char_num  ,          //字符号
    output   [511:0]   char                 //字符输出

);


always @(posedge sys_clk or negedge sys_rst_n) begin
    if(!sys_rst_n) begin
        char <= 16'd0;
    end    
    else begin
            case(char_num)
                16'd48 : char <=    512'h00000018244242424242424224180000;    //"0"
                16'd49 : char <=    512'h000000083808080808080808083E0000;    //"1"   
                16'd50 : char <=    512'h0000003C4242420204081020427E0000;    //"2"
                16'd51 : char <=    512'h0000003C4242020418040242423C0000;    //"3"
                16'd52 : char <=    512'h000000040C0C142424447F04041F0000;    //"4"
                16'd53 : char <=    512'h0000007E404040784402024244380000;    //"5"
                16'd54 : char <=    512'h000000182440405C62424242221C0000;    //"6"   
                16'd55 : char <=    512'h0000007E420404080810101010100000;    //"7"
                16'd56 : char <=    512'h0000003C4242422418244242423C0000;    //"8"
                16'd57 : char <=    512'h0000003844424242463A020224180000;    //"9"
                default : char <=   512'h00000000000000000000000000000000;
            endcase    
    end
end    


endmodule
